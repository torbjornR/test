Entety blaha.
port(

    );
